    ����          Assembly-CSharp   PauseGame+PlayerSave   xyzCHPMaxHP        ���~�aB   �  �B  �B