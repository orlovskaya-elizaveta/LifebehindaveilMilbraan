    ����          Assembly-CSharp   PauseGame+PlayerSave   xyzCHPMaxHP        �o�%sB   �  HB  �B